module memory (addr,write,read,data,clk);
input wire [4:0] addr;
input wire [7:0] data;
input wire read;
input wire clk;
input wire write;




endmodule